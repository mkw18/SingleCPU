library verilog;
use verilog.vl_types.all;
entity freq_vlg_check_tst is
    port(
        OCLK            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end freq_vlg_check_tst;
