library verilog;
use verilog.vl_types.all;
entity InstrROM_test is
end InstrROM_test;
