library verilog;
use verilog.vl_types.all;
entity regFile_test is
end regFile_test;
