library verilog;
use verilog.vl_types.all;
entity aluCtl_test is
end aluCtl_test;
