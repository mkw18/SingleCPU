library verilog;
use verilog.vl_types.all;
entity imm_PC_test is
end imm_PC_test;
