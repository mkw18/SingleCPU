library verilog;
use verilog.vl_types.all;
entity mux_data_vlg_vec_tst is
end mux_data_vlg_vec_tst;
