library verilog;
use verilog.vl_types.all;
entity mainCtl_test is
end mainCtl_test;
