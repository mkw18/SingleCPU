library verilog;
use verilog.vl_types.all;
entity SCPU_test is
end SCPU_test;
