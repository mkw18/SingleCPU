library verilog;
use verilog.vl_types.all;
entity mux_WriteAddr_vlg_vec_tst is
end mux_WriteAddr_vlg_vec_tst;
