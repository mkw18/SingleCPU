library verilog;
use verilog.vl_types.all;
entity mux_M2R_vlg_vec_tst is
end mux_M2R_vlg_vec_tst;
