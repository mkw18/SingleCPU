library verilog;
use verilog.vl_types.all;
entity mainCtl_vlg_vec_tst is
end mainCtl_vlg_vec_tst;
