library verilog;
use verilog.vl_types.all;
entity signExt_vlg_vec_tst is
end signExt_vlg_vec_tst;
